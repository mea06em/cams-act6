netcdf S5P_NRTI_L2__O3_____20240818T120300_20240818T120800_35484_03_020601_20240818T124850 {

// global attributes:
		:Conventions = "CF-1.7" ;
		:institution = "DLR-IMF" ;
		:source = "Sentinel 5 precursor, TROPOMI, space-borne remote sensing, L2" ;
		:history = "2024-08-18 12:49:05.739787 f_s5pops upas-l2 JobOrder.674317873.xml " ;
		:summary = "TROPOMI/S5P L2 data Swath 5.5x3.5km2 processed in NRTI mode" ;
		:tracking_id = "debfd6e9-b359-4f36-9f33-643cdb9e5b0b" ;
		:id = "S5P_NRTI_L2__O3_____20240818T120300_20240818T120800_35484_03_020601_20240818T124850" ;
		:time_reference = "2024-08-18T00:00:00Z" ;
		:time_reference_days_since_1950 = 27258 ;
		:time_reference_julian_day = 2460540.5 ;
		:time_reference_seconds_since_1970 = 1723939200LL ;
		:time_coverage_start = "2024-08-18T12:02:54Z" ;
		:time_coverage_end = "2024-08-18T12:08:07Z" ;
		:time_coverage_duration = "PT313.000S" ;
		:time_coverage_resolution = "PT0.840S" ;
		:orbit = 35484 ;
		:references = "TBD" ;
		:processor_version = "02.06.01" ;
		:keywords_vocabulary = "AGU index terms, http://publications.agu.org/author-resource-center/index-terms/" ;
		:keywords = "0325 Evolution of the atmosphere; 0340 Middle atmosphere, composition and chemistry; 0365 Troposphere, composition and chemistry; 1610 Atmosphere; 1630 Impacts of global change; 1640 Remote sensing" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast Metadata Conventions Standard Name Table (v29, 08 July 2015), http://cfconventions.org/standard-names.html" ;
		:naming_authority = "DLR-IMF" ;
		:cdm_data_type = "Swath" ;
		:date_created = "2024-08-18T12:49:05Z" ;
		:creator_name = "The Sentinel 5 Precursor TROPOMI Level 2 products are developed with funding from the European Space Agency (ESA), the Netherlands Space Office (NSO), the Belgian Science Policy Office, the German Aerospace Center (DLR) and the Bayerisches Staatsministerium für Wirtschaft und Medien, Energie und Technologie (StMWi)." ;
		:creator_url = "https://atmos.eoc.dlr.de/tropomi ; https://sentinel.esa.int/web/sentinel/missions/sentinel-5p" ;
		:creator_email = "EOSupport@Copernicus.esa.int" ;
		:project = "Sentinel 5 precursor/TROPOMI" ;
		:geospatial_lat_min = 33.83152f ;
		:geospatial_lat_max = 58.02542f ;
		:geospatial_lon_min = -11.08549f ;
		:geospatial_lon_max = 30.23926f ;
		:license = "No conditions apply" ;
		:platform = "S5P" ;
		:sensor = "TROPOMI" ;
		:spatial_resolution = "5.5x3.5km2" ;
		:cpp_compiler_version = "/usr/bin/c++ version 7.3.1 20180307 [gcc-7-branch revision 258314] (SUSE Linux)" ;
		:cpp_compiler_flags = "-std=gnu++11 -O2 -fopenmp" ;
		:f90_compiler_version = "/usr/bin/gfortran version 7.3.1 20180307 [gcc-7-branch revision 258314] (SUSE Linux)" ;
		:f90_compiler_flags = "-frecursive -Wno-aggressive-loop-optimizations -O2 -fopenmp" ;
		:exe_linker_flags = "-static-libgcc -static-libstdc++ -static-libgfortran" ;
		:build_date = "2023-11-10T14:17:48Z" ;
		:revision_control_identifier = "b00a2664f80dc489c4d29fdfd946e248b224a036" ;
		:geolocation_grid_from_band = 3 ;
		:identifier_product_doi = "N/A" ;
		:identifier_product_doi_authority = "http://dx.doi.org/" ;
		:algorithm_version = "UPAS-O3-DOAS_CAL-5.1.0" ;
		:product_version = "2.1" ;
		:processing_status = "Nominal" ;
		:cloud_mode = "cal" ;
		:title = "TROPOMI/S5P Ozone Total Column" ;
		:Status_MET_2D = "Nominal" ;
		:Status_NISE__ = "Nominal" ;
		:Status_L2__CLOUD_ = "External" ;
		:Status_reference_spectrum = "solar" ;
		:Status_BG = "Nominal" ;

group: PRODUCT {
  dimensions:
  	scanline = 357 ;
  	ground_pixel = 450 ;
  	time = 1 ;
  	corner = 4 ;
  	layer = 13 ;
  	level = 14 ;
  variables:
  	int scanline(scanline) ;
  		scanline:_FillValue = -2147483647 ;
  		scanline:units = "1" ;
  		scanline:axis = "Y" ;
  		scanline:long_name = "along-track dimension index" ;
  		scanline:comment = "This coordinate variable defines the indices along track; index starts at 0" ;
  	int ground_pixel(ground_pixel) ;
  		ground_pixel:_FillValue = -2147483647 ;
  		ground_pixel:units = "1" ;
  		ground_pixel:axis = "X" ;
  		ground_pixel:long_name = "across-track dimension index" ;
  		ground_pixel:comment = "This coordinate variable defines the indices across track, from west to east; index starts at 0" ;
  	int time(time) ;
  		time:_FillValue = -2147483647 ;
  		time:units = "seconds since 2010-01-01 00:00:00" ;
  		time:standard_name = "time" ;
  		time:axis = "T" ;
  		time:long_name = "reference time for the measurements" ;
  		time:comment = "The time in this variable corresponds to the time in the time_reference global attribute" ;
  	int corner(corner) ;
  		corner:_FillValue = -2147483647 ;
  		corner:units = "1" ;
  		corner:long_name = "pixel corner index" ;
  		corner:comment = "This coordinate variable defines the indices for the pixel corners; index starts a 0 (counter-clockwise, starting from south-western corner of the pixel in ascending part of the orbit)." ;
  	float latitude(time, scanline, ground_pixel) ;
  		latitude:_FillValue = 9.96921e+36f ;
  		latitude:long_name = "pixel center latitude" ;
  		latitude:units = "degrees_north" ;
  		latitude:standard_name = "latitude" ;
  		latitude:valid_min = -90.f ;
  		latitude:valid_max = 90.f ;
  		latitude:bounds = "/PRODUCT/SUPPORT_DATA/GEOLOCATIONS/latitude_bounds" ;
  	float longitude(time, scanline, ground_pixel) ;
  		longitude:_FillValue = 9.96921e+36f ;
  		longitude:long_name = "pixel center longitude" ;
  		longitude:units = "degrees_east" ;
  		longitude:standard_name = "longitude" ;
  		longitude:valid_min = -180.f ;
  		longitude:valid_max = 180.f ;
  		longitude:bounds = "/PRODUCT/SUPPORT_DATA/GEOLOCATIONS/longitude_bounds" ;
  	int delta_time(time, scanline, ground_pixel) ;
  		delta_time:_FillValue = -2147483647 ;
  		delta_time:long_name = "offset from reference start time of measurement" ;
  		delta_time:units = "milliseconds since 2024-08-18 00:00:00Z" ;
  	string time_utc(time, scanline) ;
  		string time_utc:_FillValue = "" ;
  		time_utc:long_name = "Time of observation as ISO 8601 date-time string" ;
  	ubyte qa_value(time, scanline, ground_pixel) ;
  		qa_value:_FillValue = 255UB ;
  		qa_value:units = "1" ;
  		qa_value:scale_factor = 0.01f ;
  		qa_value:add_offset = 0.f ;
  		qa_value:valid_min = 0UB ;
  		qa_value:valid_max = 100UB ;
  		qa_value:long_name = "data quality value" ;
  		qa_value:comment = "A continuous quality descriptor, varying between 0 (no data) and 1 (full quality data). Recommend to ignore data with qa_value < 0.5" ;
  		qa_value:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
  	float ozone_total_vertical_column(time, scanline, ground_pixel) ;
  		ozone_total_vertical_column:_FillValue = 9.96921e+36f ;
  		ozone_total_vertical_column:units = "mol m-2" ;
  		ozone_total_vertical_column:standard_name = "atmosphere_mole_content_of_ozone" ;
  		ozone_total_vertical_column:long_name = "total ozone column" ;
  		ozone_total_vertical_column:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
  		ozone_total_vertical_column:multiplication_factor_to_convert_to_DU = 2241.15f ;
  		ozone_total_vertical_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
  	float ozone_total_vertical_column_precision(time, scanline, ground_pixel) ;
  		ozone_total_vertical_column_precision:_FillValue = 9.96921e+36f ;
  		ozone_total_vertical_column_precision:units = "mol m-2" ;
  		ozone_total_vertical_column_precision:standard_name = "atmosphere_mole_content_of_ozone error" ;
  		ozone_total_vertical_column_precision:long_name = "total ozone column random error" ;
  		ozone_total_vertical_column_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
  		ozone_total_vertical_column_precision:multiplication_factor_to_convert_to_DU = 2241.15f ;
  		ozone_total_vertical_column_precision:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
  	int layer(layer) ;
  		layer:units = "1" ;
  		layer:long_name = "layer dimension index" ;
  	int level(level) ;
  		level:units = "1" ;
  		level:long_name = "level dimension index" ;

  group: SUPPORT_DATA {

    group: INPUT_DATA {
      variables:
      	float surface_altitude(time, scanline, ground_pixel) ;
      		surface_altitude:_FillValue = 9.96921e+36f ;
      		surface_altitude:long_name = "surface altitude" ;
      		surface_altitude:standard_name = "surface_altitude" ;
      		surface_altitude:units = "m" ;
      		surface_altitude:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_altitude:source = "http://topotools.cr.usgs.gov/gmted_viewer/" ;
      		surface_altitude:comment = "The mean of the sub-pixels of the surface altitude above the reference geoid (WGS84) within the approximate field of view, based on the GMTED2010 surface elevation database" ;
      	float surface_altitude_precision(time, scanline, ground_pixel) ;
      		surface_altitude_precision:_FillValue = 9.96921e+36f ;
      		surface_altitude_precision:long_name = "surface altitude precision" ;
      		surface_altitude_precision:standard_name = "surface_altitude standard_error" ;
      		surface_altitude_precision:units = "m" ;
      		surface_altitude_precision:standard_error_multiplier = 1.f ;
      		surface_altitude_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		surface_altitude_precision:source = "http://topotools.cr.usgs.gov/gmted_viewer/" ;
      		surface_altitude_precision:comment = "The standard deviation of sub-pixels used in calculating the mean surface altitude above the reference geoid (WGS84) within the approximate field of view, based on the GMTED2010 surface elevation database" ;
      	ubyte surface_classification(time, scanline, ground_pixel) ;
      		surface_classification:_FillValue = 255UB ;
      		surface_classification:units = "1" ;
      		surface_classification:long_name = "land-water mask" ;
      		surface_classification:comment = "flag indicating land/water and further surface classifications for the ground pixel" ;
      		surface_classification:source = "USGS (http://edc2.usgs.gov/glcc/globdoc2_0.php) and NASA SDP toolkit (http://newsroom.gsfc.nasa.gov/sdptoolkit/toolkit.html)" ;
      		surface_classification:flag_meanings = "land, water, some_water, coast, value_covers_majority_of_pixel, water+shallow_ocean, water+shallow_inland_water, water+ocean_coastline-lake_shoreline, water+intermittent_water, water+deep_inland_water, water+continental_shelf_ocean, water+deep_ocean, land+urban_and_built-up_land, land+dryland_cropland_and_pasture, land+irrigated_cropland_and_pasture, land+mixed_dryland-irrigated_cropland_and_pasture, land+cropland-grassland_mosaic, land+cropland-woodland_mosaic, land+grassland, land+shrubland, land+mixed_shrubland-grassland, land+savanna, land+deciduous_broadleaf_forest, land+deciduous_needleleaf_forest, land+evergreen_broadleaf_forest, land+evergreen_needleleaf_forest, land+mixed_forest, land+herbaceous_wetland, land+wooded_wetland, land+barren_or_sparsely_vegetated, land+herbaceous_tundra, land+wooded_tundra, land+mixed_tundra, land+bare_ground_tundra, land+snow_or_ice" ;
      		surface_classification:flag_values = 0UB, 1UB, 2UB, 3UB, 4UB, 9UB, 17UB, 25UB, 33UB, 41UB, 49UB, 57UB, 8UB, 16UB, 24UB, 32UB, 40UB, 48UB, 56UB, 64UB, 72UB, 80UB, 88UB, 96UB, 104UB, 112UB, 120UB, 128UB, 136UB, 144UB, 152UB, 160UB, 168UB, 176UB, 184UB ;
      		surface_classification:flag_masks = 3UB, 3UB, 3UB, 3UB, 4UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB, 249UB ;
      		surface_classification:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	int instrument_configuration_identifier(time, scanline) ;
      		instrument_configuration_identifier:_FillValue = -2147483647 ;
      		instrument_configuration_identifier:long_name = "IcID" ;
      		instrument_configuration_identifier:comment = "The Instrument Configuration ID defines the type of measurement and its purpose. The number of instrument configuration IDs will increase over the mission as new types of measurements are created and used" ;
      	short instrument_configuration_version(time, scanline) ;
      		instrument_configuration_version:_FillValue = -32767s ;
      		instrument_configuration_version:long_name = "IcVersion" ;
      		instrument_configuration_version:comment = "Version of the instrument_configuration_identifier" ;
      	float scaled_small_pixel_variance(time, scanline, ground_pixel) ;
      		scaled_small_pixel_variance:_FillValue = 9.96921e+36f ;
      		scaled_small_pixel_variance:long_name = "scaled small pixel variance" ;
      		scaled_small_pixel_variance:units = "1" ;
      		scaled_small_pixel_variance:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		scaled_small_pixel_variance:comment = "The scaled variance of the reflectances of the small pixels" ;
      		scaled_small_pixel_variance:radiation_wavelength = "" ;
      	float surface_pressure(time, scanline, ground_pixel) ;
      		surface_pressure:_FillValue = 9.96921e+36f ;
      		surface_pressure:units = "Pa" ;
      		surface_pressure:standard_name = "surface_air_pressure" ;
      		surface_pressure:long_name = "surface_air_pressure" ;
      		surface_pressure:source = "" ;
      		surface_pressure:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float surface_temperature(time, scanline, ground_pixel) ;
      		surface_temperature:_FillValue = 9.96921e+36f ;
      		surface_temperature:units = "K" ;
      		surface_temperature:standard_name = "surface_air_temperature" ;
      		surface_temperature:long_name = "surface_air_temperature" ;
      		surface_temperature:source = "" ;
      		surface_temperature:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float northward_wind(time, scanline, ground_pixel) ;
      		northward_wind:_FillValue = 9.96921e+36f ;
      		northward_wind:units = "m s-1" ;
      		northward_wind:standard_name = "northward_wind" ;
      		northward_wind:long_name = "Northward wind from ECMWF at 10 meter height level" ;
      		northward_wind:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float eastward_wind(time, scanline, ground_pixel) ;
      		eastward_wind:_FillValue = 9.96921e+36f ;
      		eastward_wind:units = "m s-1" ;
      		eastward_wind:standard_name = "eastward_wind" ;
      		eastward_wind:long_name = "Eastward wind from ECMWF at 10 meter height level" ;
      		eastward_wind:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_fraction(time, scanline, ground_pixel) ;
      		cloud_fraction:_FillValue = 9.96921e+36f ;
      		cloud_fraction:units = "1" ;
      		cloud_fraction:long_name = "effective radiometric cloud fraction" ;
      		cloud_fraction:source = "cal" ;
      		cloud_fraction:comment = "Coregistered effective radiometric cloud fraction using the OCRA/ROCINN CAL model." ;
      		cloud_fraction:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_fraction_precision(time, scanline, ground_pixel) ;
      		cloud_fraction_precision:_FillValue = 9.96921e+36f ;
      		cloud_fraction_precision:units = "1" ;
      		cloud_fraction_precision:long_name = "effective radiometric cloud fraction precision" ;
      		cloud_fraction_precision:source = "cal" ;
      		cloud_fraction_precision:comment = "Error of the coregistered effective radiometric cloud fraction using the OCRA/ROCINN CAL model." ;
      		cloud_fraction_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_top_pressure(time, scanline, ground_pixel) ;
      		cloud_top_pressure:_FillValue = 9.96921e+36f ;
      		cloud_top_pressure:units = "Pa" ;
      		cloud_top_pressure:standard_name = "air_pressure_at_cloud_top" ;
      		cloud_top_pressure:long_name = "cloud optical centroid top pressure" ;
      		cloud_top_pressure:source = "cal" ;
      		cloud_top_pressure:comment = "Coregistered and converted atmospheric pressure at the level of cloud top using the OCRA/ROCINN CAL model." ;
      		cloud_top_pressure:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_top_pressure_precision(time, scanline, ground_pixel) ;
      		cloud_top_pressure_precision:_FillValue = 9.96921e+36f ;
      		cloud_top_pressure_precision:units = "Pa" ;
      		cloud_top_pressure_precision:standard_name = "air_pressure_at_cloud_top standard_error" ;
      		cloud_top_pressure_precision:long_name = "cloud optical centroid top pressure precision" ;
      		cloud_top_pressure_precision:source = "cal" ;
      		cloud_top_pressure_precision:comment = "Error of the coregistered and converted atmospheric pressure at the level of cloud top using the OCRA/ROCINN CAL model." ;
      		cloud_top_pressure_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_base_pressure(time, scanline, ground_pixel) ;
      		cloud_base_pressure:_FillValue = 9.96921e+36f ;
      		cloud_base_pressure:units = "Pa" ;
      		cloud_base_pressure:standard_name = "air_pressure_at_cloud_base" ;
      		cloud_base_pressure:long_name = "cloud base pressure assumed in ROCINN retrieval" ;
      		cloud_base_pressure:source = "cal" ;
      		cloud_base_pressure:comment = "Coregistered and converted cloud base pressure retrieved using the OCRA/ROCINN CAL model." ;
      		cloud_base_pressure:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_base_pressure_precision(time, scanline, ground_pixel) ;
      		cloud_base_pressure_precision:_FillValue = 9.96921e+36f ;
      		cloud_base_pressure_precision:units = "Pa" ;
      		cloud_base_pressure_precision:standard_name = "air_pressure_at_cloud_base standard_error" ;
      		cloud_base_pressure_precision:long_name = "cloud base pressure precision assumed in ROCINN retrieval" ;
      		cloud_base_pressure_precision:source = "cal" ;
      		cloud_base_pressure_precision:comment = "Error of the coregistered and converted cloud base pressure retrieved using the OCRA/ROCINN CAL model" ;
      		cloud_base_pressure_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_top_height(time, scanline, ground_pixel) ;
      		cloud_top_height:_FillValue = 9.96921e+36f ;
      		cloud_top_height:units = "m" ;
      		cloud_top_height:long_name = "cloud top height" ;
      		cloud_top_height:source = "cal" ;
      		cloud_top_height:comment = "Coregistered vertical distance of the cloud top above the surface w.r.t. the geoid/MSL using the OCRA/ROCINN CAL model." ;
      		cloud_top_height:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_top_height_precision(time, scanline, ground_pixel) ;
      		cloud_top_height_precision:_FillValue = 9.96921e+36f ;
      		cloud_top_height_precision:units = "m" ;
      		cloud_top_height_precision:long_name = "cloud top height precision" ;
      		cloud_top_height_precision:source = "cal" ;
      		cloud_top_height_precision:comment = "Error of the coregistered vertical distance of the cloud top above the surface w.r.t. the geoid/MSL using the OCRA/ROCINN CAL model." ;
      		cloud_top_height_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_base_height(time, scanline, ground_pixel) ;
      		cloud_base_height:_FillValue = 9.96921e+36f ;
      		cloud_base_height:units = "m" ;
      		cloud_base_height:long_name = "cloud base height assumed in ROCINN retrieval" ;
      		cloud_base_height:source = "cal" ;
      		cloud_base_height:comment = "Coregistered cloud base height w.r.t. the geoid/MSL using the OCRA/ROCINN CAL model." ;
      		cloud_base_height:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_base_height_precision(time, scanline, ground_pixel) ;
      		cloud_base_height_precision:_FillValue = 9.96921e+36f ;
      		cloud_base_height_precision:units = "m" ;
      		cloud_base_height_precision:long_name = "cloud base height precision assumed in ROCINN retrieval" ;
      		cloud_base_height_precision:source = "cal" ;
      		cloud_base_height_precision:comment = "Error of the coregistered cloud base height w.r.t. the geoid/MSL using the OCRA/ROCINN CAL model." ;
      		cloud_base_height_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_optical_thickness(time, scanline, ground_pixel) ;
      		cloud_optical_thickness:_FillValue = 9.96921e+36f ;
      		cloud_optical_thickness:units = "1" ;
      		cloud_optical_thickness:standard_name = "atmosphere_optical_thickness_due_to_cloud" ;
      		cloud_optical_thickness:long_name = "cloud optical thickness" ;
      		cloud_optical_thickness:source = "cal" ;
      		cloud_optical_thickness:comment = "Coregistered cloud optical thickness based on the OCRA/ROCINN CAL model." ;
      		cloud_optical_thickness:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_optical_thickness_precision(time, scanline, ground_pixel) ;
      		cloud_optical_thickness_precision:_FillValue = 9.96921e+36f ;
      		cloud_optical_thickness_precision:units = "1" ;
      		cloud_optical_thickness_precision:standard_name = "atmosphere_optical_thickness_due_to_cloud standard_error" ;
      		cloud_optical_thickness_precision:long_name = "cloud optical thickness precision coregistered using the OCRA/ROCINN CAL model." ;
      		cloud_optical_thickness_precision:source = "cal" ;
      		cloud_optical_thickness_precision:comment = "Error of the coregistered cloud optical thickness based on the OCRA/ROCINN CAL model." ;
      		cloud_optical_thickness_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	ubyte snow_ice_flag_nise(time, scanline, ground_pixel) ;
      		snow_ice_flag_nise:units = "1" ;
      		snow_ice_flag_nise:long_name = "snow-ice mask" ;
      		snow_ice_flag_nise:_FillValue = 254UB ;
      		snow_ice_flag_nise:comment = "flag indicating snow/ice at center of ground pixel" ;
      		snow_ice_flag_nise:source = "NSIDC/NISE" ;
      		snow_ice_flag_nise:flag_meanings = "snow-free_land sea_ice_1_percent sea_ice_2_percent sea_ice_3_percent sea_ice_4_percent sea_ice_5_percent sea_ice_6_percent sea_ice_7_percent sea_ice_8_percent sea_ice_9_percent sea_ice_10_percent sea_ice_11_percent sea_ice_12_percent sea_ice_13_percent sea_ice_14_percent sea_ice_15_percent sea_ice_16_percent sea_ice_17_percent sea_ice_18_percent sea_ice_19_percent sea_ice_20_percent sea_ice_21_percent sea_ice_22_percent sea_ice_23_percent sea_ice_24_percent sea_ice_25_percent sea_ice_26_percent sea_ice_27_percent sea_ice_28_percent sea_ice_29_percent sea_ice_30_percent sea_ice_31_percent sea_ice_32_percent sea_ice_33_percent sea_ice_34_percent sea_ice_35_percent sea_ice_36_percent sea_ice_37_percent sea_ice_38_percent sea_ice_39_percent sea_ice_40_percent sea_ice_41_percent sea_ice_42_percent sea_ice_43_percent sea_ice_44_percent sea_ice_45_percent sea_ice_46_percent sea_ice_47_percent sea_ice_48_percent sea_ice_49_percent sea_ice_50_percent sea_ice_51_percent sea_ice_52_percent sea_ice_53_percent sea_ice_54_percent sea_ice_55_percent sea_ice_56_percent sea_ice_57_percent sea_ice_58_percent sea_ice_59_percent sea_ice_60_percent sea_ice_61_percent sea_ice_62_percent sea_ice_63_percent sea_ice_64_percent sea_ice_65_percent sea_ice_66_percent sea_ice_67_percent sea_ice_68_percent sea_ice_69_percent sea_ice_70_percent sea_ice_71_percent sea_ice_72_percent sea_ice_73_percent sea_ice_74_percent sea_ice_75_percent sea_ice_76_percent sea_ice_77_percent sea_ice_78_percent sea_ice_79_percent sea_ice_80_percent sea_ice_81_percent sea_ice_82_percent sea_ice_83_percent sea_ice_84_percent sea_ice_85_percent sea_ice_86_percent sea_ice_87_percent sea_ice_88_percent sea_ice_89_percent sea_ice_90_percent sea_ice_91_percent sea_ice_92_percent sea_ice_93_percent sea_ice_94_percent sea_ice_95_percent sea_ice_96_percent sea_ice_97_percent sea_ice_98_percent sea_ice_99_percent sea_ice_100_percent permanent_ice snow mixed_pixels_at_coastlines suspect_ice_value corners ocean" ;
      		snow_ice_flag_nise:flag_values = 0UB, 1UB, 2UB, 3UB, 4UB, 5UB, 6UB, 7UB, 8UB, 9UB, 10UB, 11UB, 12UB, 13UB, 14UB, 15UB, 16UB, 17UB, 18UB, 19UB, 20UB, 21UB, 22UB, 23UB, 24UB, 25UB, 26UB, 27UB, 28UB, 29UB, 30UB, 31UB, 32UB, 33UB, 34UB, 35UB, 36UB, 37UB, 38UB, 39UB, 40UB, 41UB, 42UB, 43UB, 44UB, 45UB, 46UB, 47UB, 48UB, 49UB, 50UB, 51UB, 52UB, 53UB, 54UB, 55UB, 56UB, 57UB, 58UB, 59UB, 60UB, 61UB, 62UB, 63UB, 64UB, 65UB, 66UB, 67UB, 68UB, 69UB, 70UB, 71UB, 72UB, 73UB, 74UB, 75UB, 76UB, 77UB, 78UB, 79UB, 80UB, 81UB, 82UB, 83UB, 84UB, 85UB, 86UB, 87UB, 88UB, 89UB, 90UB, 91UB, 92UB, 93UB, 94UB, 95UB, 96UB, 97UB, 98UB, 99UB, 100UB, 101UB, 103UB, 252UB, 253UB, 254UB, 255UB ;
      		snow_ice_flag_nise:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	ubyte snow_ice_flag(time, scanline, ground_pixel) ;
      		snow_ice_flag:units = "1" ;
      		snow_ice_flag:threshold = "0.3" ;
      		snow_ice_flag:long_name = "snow-ice mask" ;
      		snow_ice_flag:_FillValue = 254UB ;
      		snow_ice_flag:comment = "flag indicating snow/ice at center of ground pixel" ;
      		snow_ice_flag:source = "" ;
      		snow_ice_flag:flag_meanings = "snow_free snow_ice" ;
      		snow_ice_flag:flag_values = 0UB, 1UB ;
      		snow_ice_flag:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float snow_cover(time, scanline, ground_pixel) ;
      		snow_cover:_FillValue = 9.96921e+36f ;
      		snow_cover:units = "1" ;
      		snow_cover:long_name = "snow-cover" ;
      		snow_cover:source = "ECMWF" ;
      		snow_cover:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float sea_ice_cover(time, scanline, ground_pixel) ;
      		sea_ice_cover:_FillValue = 9.96921e+36f ;
      		sea_ice_cover:units = "1" ;
      		sea_ice_cover:long_name = "sea-ice-cover" ;
      		sea_ice_cover:source = "ECMWF" ;
      		sea_ice_cover:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float surface_albedo(time, scanline, ground_pixel) ;
      		surface_albedo:_FillValue = 9.96921e+36f ;
      		surface_albedo:units = "1" ;
      		surface_albedo:standard_name = "surface_albedo" ;
      		surface_albedo:long_name = "surface albedo from daily G3_LER" ;
      		surface_albedo:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float effective_scene_height(time, scanline, ground_pixel) ;
      		effective_scene_height:_FillValue = 9.96921e+36f ;
      		effective_scene_height:units = "m" ;
      		effective_scene_height:standard_name = "TBD" ;
      		effective_scene_height:long_name = "effective scene height from the CRB model" ;
      		effective_scene_height:source = "crb" ;
      		effective_scene_height:comment = "Effective Scene Height using the OCRA/ROCINN CRB model." ;
      		effective_scene_height:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float effective_scene_height_precision(time, scanline, ground_pixel) ;
      		effective_scene_height_precision:_FillValue = 9.96921e+36f ;
      		effective_scene_height_precision:units = "m" ;
      		effective_scene_height_precision:standard_name = "TBD" ;
      		effective_scene_height_precision:long_name = "effective scene height precision from the CRB model" ;
      		effective_scene_height_precision:source = "crb" ;
      		effective_scene_height_precision:comment = "Error of the effective scene height using the OCRA/ROCINN CRB model." ;
      		effective_scene_height_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float effective_scene_pressure(time, scanline, ground_pixel) ;
      		effective_scene_pressure:_FillValue = 9.96921e+36f ;
      		effective_scene_pressure:units = "Pa" ;
      		effective_scene_pressure:standard_name = "TBD" ;
      		effective_scene_pressure:long_name = "effective scene optical centroid pressure from the CRB model" ;
      		effective_scene_pressure:source = "crb" ;
      		effective_scene_pressure:comment = "Effective scene pressure using the OCRA/ROCINN CRB model." ;
      		effective_scene_pressure:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float effective_scene_pressure_precision(time, scanline, ground_pixel) ;
      		effective_scene_pressure_precision:_FillValue = 9.96921e+36f ;
      		effective_scene_pressure_precision:units = "Pa" ;
      		effective_scene_pressure_precision:standard_name = "TBD" ;
      		effective_scene_pressure_precision:long_name = "effective scene pressure precision from the CRB model" ;
      		effective_scene_pressure_precision:source = "crb" ;
      		effective_scene_pressure_precision:comment = "Error of the effective scene pressure using the OCRA/ROCINN CRB model." ;
      		effective_scene_pressure_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_fraction_apriori(time, scanline, ground_pixel) ;
      		cloud_fraction_apriori:_FillValue = 9.96921e+36f ;
      		cloud_fraction_apriori:units = "1" ;
      		cloud_fraction_apriori:long_name = "effective radiometric cloud fraction a priori" ;
      		cloud_fraction_apriori:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;

      group: PROCESSOR {

        // group attributes:
        		:processing_configuration = "./upas-l2 --time-slot 20240818T120300.000000-20240818T120800.000000 -d /mnt/sw/IPF_S5P_L2_DLR/current/processors/support_data -t 26 -m NRTI --degradation-step-acrosstrack 0 --degradation-step-alongtrack 0 -e 2024-08-18 12:49:05.739787 f_s5pops upas-l2 JobOrder.674317873.xml PDGS-OP --o3 -o /mnt/data1/storage_nrt/cache_nrt/O3-674319189/S5P_NRTI_L2__O3_____20240818T120300_20240818T120800_35484_03_020601_20240818T124850.nc /mnt/data1/storage_nrt/cache_nrt/AUX_O3-674319170/S5P_OFFL_L1B_IR_UVN_20240817T162923_20240817T181053_35473_03_020100_20240818T030032.nc /mnt/data1/storage_nrt/cache_nrt/L1B-674317875/S5P_NRTI_L1B_RA_BD1_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc /mnt/data1/storage_nrt/cache_nrt/L1B-674317875/S5P_NRTI_L1B_RA_BD2_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc /mnt/data1/storage_nrt/cache_nrt/L1B-674317875/S5P_NRTI_L1B_RA_BD3_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc /mnt/data1/storage_nrt/cache_nrt/L1B-674317875/S5P_NRTI_L1B_RA_BD4_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc /mnt/data1/storage_nrt/cache_nrt/L1B-674317875/S5P_NRTI_L1B_RA_BD5_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc /mnt/data1/storage_nrt/cache_nrt/L1B-674317875/S5P_NRTI_L1B_RA_BD6_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc /mnt/data1/storage_nrt/cache_nrt/L1B-674317875/S5P_NRTI_L1B_RA_BD7_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc /mnt/data1/storage_nrt/cache_nrt/L1B-674317875/S5P_NRTI_L1B_RA_BD8_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc --aux-cloud /mnt/data1/storage_nrt/cache_nrt/CLOUD-674319180/S5P_NRTI_L2__CLOUD__20240818T120300_20240818T120800_35484_03_020601_20240818T124206.nc --aux-bgo3 /mnt/data1/storage_nrt/pp_bgo3/S5P_NRTI_AUX_BGO3___20240815T205808_20240817T000320_20240818T000018.nc " ;
        } // group PROCESSOR
      } // group INPUT_DATA

    group: GEOLOCATIONS {
      variables:
      	float satellite_latitude(time, scanline) ;
      		satellite_latitude:_FillValue = 9.96921e+36f ;
      		satellite_latitude:long_name = "sub satellite latitude" ;
      		satellite_latitude:units = "degrees_north" ;
      		satellite_latitude:comment = "Latitude of the geodetic sub satellite point on the WGS84 reference ellipsoid" ;
      		satellite_latitude:valid_min = -90.f ;
      		satellite_latitude:valid_max = 90.f ;
      	float satellite_longitude(time, scanline) ;
      		satellite_longitude:_FillValue = 9.96921e+36f ;
      		satellite_longitude:long_name = "satellite_longitude" ;
      		satellite_longitude:units = "degrees_east" ;
      		satellite_longitude:comment = "Longitude of the geodetic sub satellite point on the WGS84 reference ellipsoid" ;
      		satellite_longitude:valid_min = -180.f ;
      		satellite_longitude:valid_max = 180.f ;
      	float satellite_altitude(time, scanline) ;
      		satellite_altitude:_FillValue = 9.96921e+36f ;
      		satellite_altitude:long_name = "satellite altitude" ;
      		satellite_altitude:units = "m" ;
      		satellite_altitude:comment = "The altitude of the satellite with respect to the geodetic sub satellite point on the WGS84 reference ellipsoid" ;
      		satellite_altitude:valid_min = 700000.f ;
      		satellite_altitude:valid_max = 900000.f ;
      	float satellite_orbit_phase(time, scanline) ;
      		satellite_orbit_phase:_FillValue = 9.96921e+36f ;
      		satellite_orbit_phase:long_name = "fractional satellite orbit phase" ;
      		satellite_orbit_phase:units = "1" ;
      		satellite_orbit_phase:comment = "Relative offset [0.0, ..., 1.0] of the measurement in the orbit" ;
      		satellite_orbit_phase:valid_min = -0.02f ;
      		satellite_orbit_phase:valid_max = 1.02f ;
      	float solar_zenith_angle(time, scanline, ground_pixel) ;
      		solar_zenith_angle:_FillValue = 9.96921e+36f ;
      		solar_zenith_angle:long_name = "solar zenith angle" ;
      		solar_zenith_angle:standard_name = "solar_zenith_angle" ;
      		solar_zenith_angle:units = "degree" ;
      		solar_zenith_angle:valid_min = 0.f ;
      		solar_zenith_angle:valid_max = 180.f ;
      		solar_zenith_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		solar_zenith_angle:comment = "Solar zenith angle at the ground pixel location on the reference ellipsoid. Angle is measured away from the vertical" ;
      	float solar_azimuth_angle(time, scanline, ground_pixel) ;
      		solar_azimuth_angle:_FillValue = 9.96921e+36f ;
      		solar_azimuth_angle:long_name = "solar azimuth angle" ;
      		solar_azimuth_angle:standard_name = "solar_azimuth_angle" ;
      		solar_azimuth_angle:units = "degree" ;
      		solar_azimuth_angle:valid_min = -180.f ;
      		solar_azimuth_angle:valid_max = 180.f ;
      		solar_azimuth_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		solar_azimuth_angle:comment = "Solar azimuth angle at the ground pixel location on the reference ellipsoid. Angle is measured clockwise from the North (East = 90, South = +/-180, West = -90)" ;
      	float viewing_zenith_angle(time, scanline, ground_pixel) ;
      		viewing_zenith_angle:_FillValue = 9.96921e+36f ;
      		viewing_zenith_angle:long_name = "viewing zenith angle" ;
      		viewing_zenith_angle:standard_name = "viewing_zenith_angle" ;
      		viewing_zenith_angle:units = "degree" ;
      		viewing_zenith_angle:valid_min = 0.f ;
      		viewing_zenith_angle:valid_max = 180.f ;
      		viewing_zenith_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		viewing_zenith_angle:comment = "Zenith angle of the satellite at the ground pixel location on the reference ellipsoid. Angle is measured away from the vertical" ;
      	float viewing_azimuth_angle(time, scanline, ground_pixel) ;
      		viewing_azimuth_angle:_FillValue = 9.96921e+36f ;
      		viewing_azimuth_angle:long_name = "viewing azimuth angle" ;
      		viewing_azimuth_angle:standard_name = "viewing_azimuth_angle" ;
      		viewing_azimuth_angle:units = "degree" ;
      		viewing_azimuth_angle:valid_min = -180.f ;
      		viewing_azimuth_angle:valid_max = 180.f ;
      		viewing_azimuth_angle:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		viewing_azimuth_angle:comment = "Satellite azimuth angle at the ground pixel location on the reference ellipsoid. Angle is measured clockwise from the North (East = 90, South = +/-180, West = -90)" ;
      	float latitude_bounds(time, scanline, ground_pixel, corner) ;
      		latitude_bounds:_FillValue = 9.96921e+36f ;
      		latitude_bounds:units = "degrees_north" ;
      	float longitude_bounds(time, scanline, ground_pixel, corner) ;
      		longitude_bounds:_FillValue = 9.96921e+36f ;
      		longitude_bounds:units = "degrees_east" ;
      	ubyte geolocation_flags(time, scanline, ground_pixel) ;
      		geolocation_flags:_FillValue = 255UB ;
      		geolocation_flags:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		geolocation_flags:flag_masks = 0UB, 1UB, 2UB, 4UB, 8UB, 16UB, 32UB, 128UB ;
      		geolocation_flags:flag_meanings = "no_error solar_eclipse sun_glint_possible descending night geo_boundary_crossing spacecraft_manoeuvre geolocation_error" ;
      		geolocation_flags:flag_values = 0UB, 1UB, 2UB, 4UB, 8UB, 16UB, 32UB, 128UB ;
      		geolocation_flags:long_name = "geolocation flags" ;
      		geolocation_flags:max_val = 254UB ;
      		geolocation_flags:min_val = 0UB ;
      		geolocation_flags:units = "1" ;
      } // group GEOLOCATIONS

    group: DETAILED_RESULTS {
      dimensions:
      	number_of_slant_columns = 4 ;
      	number_of_doas_polynomial_coefficients = 4 ;
      variables:
      	float ozone_profile_apriori(time, scanline, ground_pixel, layer) ;
      		ozone_profile_apriori:_FillValue = 9.96921e+36f ;
      		ozone_profile_apriori:units = "mol m-2" ;
      		ozone_profile_apriori:long_name = "apriori ozone profile" ;
      		ozone_profile_apriori:positive = "up" ;
      		ozone_profile_apriori:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		ozone_profile_apriori:multiplication_factor_to_convert_to_DU = 2241.15f ;
      		ozone_profile_apriori:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      	float averaging_kernel(time, scanline, ground_pixel, layer) ;
      		averaging_kernel:_FillValue = 9.96921e+36f ;
      		averaging_kernel:units = "1" ;
      		averaging_kernel:long_name = "ozone averaging kernel" ;
      		averaging_kernel:positive = "up" ;
      		averaging_kernel:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float pressure_grid(time, scanline, ground_pixel, level) ;
      		pressure_grid:_FillValue = 9.96921e+36f ;
      		pressure_grid:units = "Pa" ;
      		pressure_grid:standard_name = "atmosphere_hybrid_sigma_pressure_coordinate" ;
      		pressure_grid:long_name = "pressure grid" ;
      		pressure_grid:positive = "up" ;
      		pressure_grid:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		pressure_grid:index_meaning = "1" ;
      	double fitted_slant_columns(time, scanline, ground_pixel, number_of_slant_columns) ;
      		fitted_slant_columns:_FillValue = 9.96920996838687e+36 ;
      		fitted_slant_columns:units = "mol m-2" ;
      		fitted_slant_columns:long_name = "slant column densities" ;
      		fitted_slant_columns:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		fitted_slant_columns:index_meaning = "O3_Brion_vac_Qparam_Full_resolution_320340_243K_NOMOPS_BF2bd2-6_band_3#1#float64#2#451x399.bis O3Diff_Brion_vac_Qparam_Full_resolution_320340_243-223K_NOMOPS_BF2bd2-6_band_3.xs#1#float64#2#451x399.bis no2_VANDAELE_1998_220K_NOMOPS_BF2bd2-6_band_3.xs#1#float64#2#451x2010.bis ring_sao2010_hr_norm_NOMOPS_BF2bd2-6_band_3#1#float64#2#451x2010.bis " ;
      		fitted_slant_columns:multiplication_factor_to_convert_to_DU = 2241.15f ;
      		fitted_slant_columns:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      	float fitted_slant_columns_precision(time, scanline, ground_pixel, number_of_slant_columns) ;
      		fitted_slant_columns_precision:_FillValue = 9.96921e+36f ;
      		fitted_slant_columns_precision:units = "mol m-2" ;
      		fitted_slant_columns_precision:long_name = "slant column density random error" ;
      		fitted_slant_columns_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		fitted_slant_columns_precision:index_meaning = "O3_Brion_vac_Qparam_Full_resolution_320340_243K_NOMOPS_BF2bd2-6_band_3#1#float64#2#451x399.bis O3Diff_Brion_vac_Qparam_Full_resolution_320340_243-223K_NOMOPS_BF2bd2-6_band_3.xs#1#float64#2#451x399.bis no2_VANDAELE_1998_220K_NOMOPS_BF2bd2-6_band_3.xs#1#float64#2#451x2010.bis ring_sao2010_hr_norm_NOMOPS_BF2bd2-6_band_3#1#float64#2#451x2010.bis " ;
      		fitted_slant_columns_precision:multiplication_factor_to_convert_to_DU = 2241.15f ;
      		fitted_slant_columns_precision:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      	ushort number_of_iterations_slant_column(time, scanline, ground_pixel) ;
      		number_of_iterations_slant_column:_FillValue = 65535US ;
      		number_of_iterations_slant_column:units = "1" ;
      		number_of_iterations_slant_column:long_name = "number of doas fit iterations" ;
      		number_of_iterations_slant_column:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float fitted_root_mean_square(time, scanline, ground_pixel) ;
      		fitted_root_mean_square:_FillValue = 9.96921e+36f ;
      		fitted_root_mean_square:units = "1" ;
      		fitted_root_mean_square:long_name = "doas fit root mean square residual" ;
      		fitted_root_mean_square:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float fitted_radiance_shift(time, scanline, ground_pixel) ;
      		fitted_radiance_shift:_FillValue = 9.96921e+36f ;
      		fitted_radiance_shift:units = "nm" ;
      		fitted_radiance_shift:long_name = "radiance wavelength shift from the doas fit" ;
      		fitted_radiance_shift:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float fitted_radiance_squeeze(time, scanline, ground_pixel) ;
      		fitted_radiance_squeeze:_FillValue = 9.96921e+36f ;
      		fitted_radiance_squeeze:units = "1" ;
      		fitted_radiance_squeeze:long_name = "radiance wavelength squeeze/stretch from the doas fit" ;
      		fitted_radiance_squeeze:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float ozone_slant_column_ring_corrected(time, scanline, ground_pixel) ;
      		ozone_slant_column_ring_corrected:_FillValue = 9.96921e+36f ;
      		ozone_slant_column_ring_corrected:units = "mol m-2" ;
      		ozone_slant_column_ring_corrected:long_name = "ring corrected slant column" ;
      		ozone_slant_column_ring_corrected:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		ozone_slant_column_ring_corrected:multiplication_factor_to_convert_to_DU = 2241.15f ;
      		ozone_slant_column_ring_corrected:multiplication_factor_to_convert_to_molecules_percm2 = 6.02214e+19f ;
      	ushort number_of_spectral_points_in_retrieval(time, scanline, ground_pixel) ;
      		number_of_spectral_points_in_retrieval:_FillValue = 65535US ;
      		number_of_spectral_points_in_retrieval:long_name = "Number of spectral points used in the DOAS retrieval" ;
      		number_of_spectral_points_in_retrieval:units = "1" ;
      		number_of_spectral_points_in_retrieval:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float ozone_total_air_mass_factor(time, scanline, ground_pixel) ;
      		ozone_total_air_mass_factor:_FillValue = 9.96921e+36f ;
      		ozone_total_air_mass_factor:units = "1" ;
      		ozone_total_air_mass_factor:long_name = "total air mass factor" ;
      		ozone_total_air_mass_factor:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float ozone_total_air_mass_factor_trueness(time, scanline, ground_pixel) ;
      		ozone_total_air_mass_factor_trueness:_FillValue = 9.96921e+36f ;
      		ozone_total_air_mass_factor_trueness:units = "1" ;
      		ozone_total_air_mass_factor_trueness:long_name = "total air mass factor systematic error" ;
      		ozone_total_air_mass_factor_trueness:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float ozone_clear_air_mass_factor(time, scanline, ground_pixel) ;
      		ozone_clear_air_mass_factor:_FillValue = 9.96921e+36f ;
      		ozone_clear_air_mass_factor:units = "1" ;
      		ozone_clear_air_mass_factor:long_name = "cloud free air mass factor" ;
      		ozone_clear_air_mass_factor:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float ozone_clear_air_mass_factor_trueness(time, scanline, ground_pixel) ;
      		ozone_clear_air_mass_factor_trueness:_FillValue = 9.96921e+36f ;
      		ozone_clear_air_mass_factor_trueness:units = "1" ;
      		ozone_clear_air_mass_factor_trueness:long_name = "cloud free air mass factor systematic error" ;
      		ozone_clear_air_mass_factor_trueness:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float ozone_cloudy_air_mass_factor(time, scanline, ground_pixel) ;
      		ozone_cloudy_air_mass_factor:_FillValue = 9.96921e+36f ;
      		ozone_cloudy_air_mass_factor:units = "1" ;
      		ozone_cloudy_air_mass_factor:long_name = "cloudy air mass factor" ;
      		ozone_cloudy_air_mass_factor:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float ozone_cloudy_air_mass_factor_trueness(time, scanline, ground_pixel) ;
      		ozone_cloudy_air_mass_factor_trueness:_FillValue = 9.96921e+36f ;
      		ozone_cloudy_air_mass_factor_trueness:units = "1" ;
      		ozone_cloudy_air_mass_factor_trueness:long_name = "cloudy air mass factor systematic error" ;
      		ozone_cloudy_air_mass_factor_trueness:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float cloud_fraction_intensity_weighted(time, scanline, ground_pixel) ;
      		cloud_fraction_intensity_weighted:_FillValue = 9.96921e+36f ;
      		cloud_fraction_intensity_weighted:units = "1" ;
      		cloud_fraction_intensity_weighted:long_name = "intensity weighted cloud fraction used for total amf calculation" ;
      		cloud_fraction_intensity_weighted:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float ozone_effective_temperature(time, scanline, ground_pixel) ;
      		ozone_effective_temperature:_FillValue = 9.96921e+36f ;
      		ozone_effective_temperature:units = "K" ;
      		ozone_effective_temperature:long_name = "ozone cross section effective temperature" ;
      		ozone_effective_temperature:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	ushort number_of_iterations_vertical_column(time, scanline, ground_pixel) ;
      		number_of_iterations_vertical_column:_FillValue = 65535US ;
      		number_of_iterations_vertical_column:units = "1" ;
      		number_of_iterations_vertical_column:long_name = "number of vcd iterations" ;
      		number_of_iterations_vertical_column:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	float effective_scene_albedo(time, scanline, ground_pixel) ;
      		effective_scene_albedo:_FillValue = 9.96921e+36f ;
      		effective_scene_albedo:units = "1" ;
      		effective_scene_albedo:long_name = "Geometry-dependent effective Lambertian equivalent reflectivity (GE_LER)" ;
      		effective_scene_albedo:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		effective_scene_albedo:comment = "GE_LER retrieved using FP_ILM" ;
      	float effective_scene_albedo_precision(time, scanline, ground_pixel) ;
      		effective_scene_albedo_precision:_FillValue = 9.96921e+36f ;
      		effective_scene_albedo_precision:units = "1" ;
      		effective_scene_albedo_precision:long_name = "GE_LER error" ;
      		effective_scene_albedo_precision:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		effective_scene_albedo_precision:comment = "Error of the GE_LER retrieved using FP_ILM" ;
      	float doas_polynomial_coefficients(time, scanline, ground_pixel, number_of_doas_polynomial_coefficients) ;
      		doas_polynomial_coefficients:_FillValue = 9.96921e+36f ;
      		doas_polynomial_coefficients:units = "1" ;
      		doas_polynomial_coefficients:long_name = "DOAS polynomial coefficients" ;
      		doas_polynomial_coefficients:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		doas_polynomial_coefficients:comment = "Values of the DOAS polynomial coefficients" ;
      	float euv(time, scanline, ground_pixel) ;
      		euv:_FillValue = 9.96921e+36f ;
      		euv:units = "W m-2" ;
      		euv:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      		euv:long_name = "Erythemal UV irradiance" ;
      	uint processing_quality_flags(time, scanline, ground_pixel) ;
      		processing_quality_flags:_FillValue = 4294967295U ;
      		processing_quality_flags:long_name = "Processing quality flags" ;
      		processing_quality_flags:units = "1" ;
      		processing_quality_flags:comment = "Flags indicating conditions that affect quality of the retrieval." ;
      		processing_quality_flags:flag_meanings = "success radiance_missing irradiance_missing input_spectrum_missing reflectance_range_error ler_range_error snr_range_error sza_range_error vza_range_error lut_range_error ozone_range_error wavelength_offset_error initialization_error memory_error assertion_error io_error numerical_error lut_error ISRF_error convergence_error cloud_filter_convergence_error max_iteration_convergence_error aot_lower_boundary_convergence_error other_boundary_convergence_error geolocation_error ch4_noscat_zero_error h2o_noscat_zero_error max_optical_thickness_error aerosol_boundary_error boundary_hit_error chi2_error svd_error dfs_error radiative_transfer_error optimal_estimation_error profile_error cloud_error model_error number_of_input_data_points_too_low_error cloud_pressure_spread_too_low_error cloud_too_low_level_error generic_range_error generic_exception input_spectrum_alignment_error abort_error wrong_input_type_error wavelength_calibration_error coregistration_error slant_column_density_error airmass_factor_error vertical_column_density_error signal_to_noise_ratio_error configuration_error key_error saturation_error max_num_outlier_exceeded_error solar_eclipse_filter cloud_filter altitude_consistency_filter altitude_roughness_filter sun_glint_filter mixed_surface_type_filter snow_ice_filter aai_filter cloud_fraction_fresco_filter aai_scene_albedo_filter small_pixel_radiance_std_filter cloud_fraction_viirs_filter cirrus_reflectance_viirs_filter cf_viirs_swir_ifov_filter cf_viirs_swir_ofova_filter cf_viirs_swir_ofovb_filter cf_viirs_swir_ofovc_filter cf_viirs_nir_ifov_filter cf_viirs_nir_ofova_filter cf_viirs_nir_ofovb_filter cf_viirs_nir_ofovc_filter refl_cirrus_viirs_swir_filter refl_cirrus_viirs_nir_filter diff_refl_cirrus_viirs_filter ch4_noscat_ratio_filter ch4_noscat_ratio_std_filter h2o_noscat_ratio_filter h2o_noscat_ratio_std_filter diff_psurf_fresco_ecmwf_filter psurf_fresco_stdv_filter ocean_filter time_range_filter pixel_or_scanline_index_filter geographic_region_filter input_spectrum_warning wavelength_calibration_warning extrapolation_warning sun_glint_warning south_atlantic_anomaly_warning sun_glint_correction snow_ice_warning cloud_warning AAI_warning pixel_level_input_data_missing data_range_warning low_cloud_fraction_warning altitude_consistency_warning signal_to_noise_ratio_warning deconvolution_warning so2_volcanic_origin_likely_warning so2_volcanic_origin_certain_warning interpolation_warning saturation_warning high_sza_warning cloud_retrieval_warning cloud_inhomogeneity_warning thermal_instability_warning" ;
      		processing_quality_flags:flag_masks = 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 255U, 256U, 512U, 1024U, 2048U, 4096U, 8192U, 16384U, 32768U, 65536U, 131072U, 262144U, 524288U, 1048576U, 2097152U, 4194304U, 8388608U, 16777216U, 33554432U, 67108864U, 134217728U, 268435456U, 536870912U, 1073741824U ;
      		processing_quality_flags:flag_values = 0U, 1U, 2U, 3U, 4U, 5U, 6U, 7U, 8U, 9U, 10U, 11U, 12U, 13U, 14U, 15U, 16U, 17U, 18U, 19U, 20U, 21U, 22U, 23U, 24U, 25U, 26U, 27U, 28U, 29U, 30U, 31U, 32U, 33U, 34U, 35U, 36U, 37U, 38U, 39U, 40U, 41U, 42U, 43U, 44U, 45U, 46U, 47U, 48U, 49U, 50U, 51U, 52U, 53U, 54U, 55U, 64U, 65U, 66U, 67U, 68U, 69U, 70U, 71U, 72U, 73U, 74U, 75U, 76U, 77U, 78U, 79U, 80U, 81U, 82U, 83U, 84U, 85U, 86U, 87U, 88U, 89U, 90U, 91U, 92U, 93U, 94U, 95U, 96U, 97U, 256U, 512U, 1024U, 2048U, 4096U, 8192U, 16384U, 32768U, 65536U, 131072U, 262144U, 524288U, 1048576U, 2097152U, 4194304U, 8388608U, 16777216U, 33554432U, 67108864U, 134217728U, 268435456U, 536870912U, 1073741824U ;
      		processing_quality_flags:coordinates = "/PRODUCT/longitude /PRODUCT/latitude" ;
      	int number_of_slant_columns(number_of_slant_columns) ;
      		number_of_slant_columns:units = "1" ;
      		number_of_slant_columns:long_name = "number_of_slant_columns dimension index" ;
      	int number_of_doas_polynomial_coefficients(number_of_doas_polynomial_coefficients) ;
      		number_of_doas_polynomial_coefficients:units = "1" ;
      		number_of_doas_polynomial_coefficients:long_name = "number_of_doas_polynomial_coefficients dimension index" ;

      group: WAVELENGTH_CALIBRATIONS {
        dimensions:
        	number_of_calibrations = 450 ;
        	degrees_of_polynomial_shift = 4 ;
        	number_of_subwindows = 4 ;
        variables:
        	float calibration_polynomial_coefficients(number_of_calibrations, degrees_of_polynomial_shift) ;
        		calibration_polynomial_coefficients:_FillValue = 9.96921e+36f ;
        		calibration_polynomial_coefficients:units = "1" ;
        		calibration_polynomial_coefficients:long_name = "computed coefficients of the polynomial function" ;
        		calibration_polynomial_coefficients:standard_name = "TBA" ;
        	float calibration_subwindows_shift(number_of_calibrations, number_of_subwindows) ;
        		calibration_subwindows_shift:_FillValue = 9.96921e+36f ;
        		calibration_subwindows_shift:units = "nm" ;
        		calibration_subwindows_shift:long_name = "irradiance wavelengths shift fitted values per subwindow" ;
        		calibration_subwindows_shift:standard_name = "TBA" ;
        	float calibration_subwindows_squeeze(number_of_calibrations, number_of_subwindows) ;
        		calibration_subwindows_squeeze:_FillValue = 9.96921e+36f ;
        		calibration_subwindows_squeeze:units = "1" ;
        		calibration_subwindows_squeeze:long_name = "irradiance wavelengths squeeze fitted values per subwindow" ;
        		calibration_subwindows_squeeze:standard_name = "TBA" ;
        	float calibration_subwindows_root_mean_square(number_of_calibrations, number_of_subwindows) ;
        		calibration_subwindows_root_mean_square:_FillValue = 9.96921e+36f ;
        		calibration_subwindows_root_mean_square:units = "1" ;
        		calibration_subwindows_root_mean_square:long_name = "calibration rms per subwindow" ;
        		calibration_subwindows_root_mean_square:standard_name = "TBA" ;
        	float calibration_subwindows_wavelength(number_of_subwindows) ;
        		calibration_subwindows_wavelength:_FillValue = 9.96921e+36f ;
        		calibration_subwindows_wavelength:units = "nm" ;
        		calibration_subwindows_wavelength:long_name = "calibration wavelength center in each subwindow" ;
        		calibration_subwindows_wavelength:standard_name = "TBA" ;
        	int number_of_calibrations(number_of_calibrations) ;
        		number_of_calibrations:units = "1" ;
        		number_of_calibrations:long_name = "number_of_calibrations dimension index" ;
        	int degrees_of_polynomial_shift(degrees_of_polynomial_shift) ;
        		degrees_of_polynomial_shift:units = "1" ;
        		degrees_of_polynomial_shift:long_name = "degrees_of_polynomial_shift dimension index" ;
        	int number_of_subwindows(number_of_subwindows) ;
        		number_of_subwindows:units = "1" ;
        		number_of_subwindows:long_name = "number_of_subwindows dimension index" ;
        } // group WAVELENGTH_CALIBRATIONS
      } // group DETAILED_RESULTS
    } // group SUPPORT_DATA
  } // group PRODUCT

group: METADATA {

  group: EOP_METADATA {

    // group attributes:
    		:gml\:id = "S5P_NRTI_L2__O3_____20240818T120300_20240818T120800_35484_03_020601_20240818T124850.ID" ;
    		:objectType = "atm:EarthObservation" ;

    group: om\:procedure {

      // group attributes:
      		:gml\:id = "S5P_NRTI_L2__O3_____20240818T120300_20240818T120800_35484_03_020601_20240818T124850.EOE" ;
      		:objectType = "eop:EarthObservationEquipment" ;

      group: eop\:sensor {

        // group attributes:
        		:eop\:sensorType = "ATMOSPHERIC" ;
        		:objectType = "eop:Sensor" ;
        } // group eop\:sensor

      group: eop\:platform {

        // group attributes:
        		:eop\:shortName = "Sentinel-5p" ;
        		:objectType = "eop:Platform" ;
        } // group eop\:platform

      group: eop\:instrument {

        // group attributes:
        		:eop\:shortName = "TROPOMI" ;
        		:objectType = "eop:Instrument" ;
        } // group eop\:instrument

      group: eop\:acquisitionParameters {

        // group attributes:
        		:eop\:orbitNumber = 35484 ;
        		:objectType = "eop:Acquisition" ;
        } // group eop\:acquisitionParameters
      } // group om\:procedure

    group: om\:phenomenonTime {

      // group attributes:
      		:gml\:beginPosition = "2024-08-18T12:02:54Z" ;
      		:gml\:endPosition = "2024-08-18T12:08:07Z" ;
      		:objectType = "gml:TimePeriod" ;
      } // group om\:phenomenonTime

    group: om\:observedProperty {

      // group attributes:
      		:nilReason = "inapplicable" ;
      } // group om\:observedProperty

    group: om\:featureOfInterest {

      // group attributes:
      		:objectType = "eop:FootPrint" ;
      		:gml\:id = "S5P_NRTI_L2__O3_____20240818T120300_20240818T120800_35484_03_020601_20240818T124850.FP" ;

      group: eop\:multiExtentOf {

        // group attributes:
        		:objectType = "gml:MultiSurface" ;

        group: gml\:surfaceMembers {

          // group attributes:
          		:objectType = "gml:Polygon" ;

          group: gml\:exterior {

            // group attributes:
            		:gml\:posList = "50.47874 -11.085491 49.203228 -9.836398 47.913067 -8.655639 46.60939 -7.5380745 45.29375 -6.4783893 43.966778 -5.472516 42.629475 -4.516469 41.282864 -3.6060276 39.927567 -2.738356 38.564404 -1.9098043 37.19383 -1.1182761 35.81647 -0.3608863 34.432922 0.36501244 33.83152 0.670182 33.87532 0.7582091 34.66445 2.3853943 35.8854 5.096727 36.599663 6.8403926 37.19815 8.439581 37.60267 9.623783 37.975193 10.818784 38.245853 11.772063 38.509846 12.794526 38.711193 13.655172 38.89948 14.543856 38.915623 14.624658 39.076725 15.479885 39.244198 16.488998 39.377914 17.42238 39.51662 18.580502 39.624676 19.71207 39.72935 21.207481 39.79794 22.782463 39.83296 25.078274 39.79024 27.853357 39.69093 30.239256 41.136562 30.100107 42.581497 29.970097 44.025723 29.84986 45.46904 29.740007 46.911564 29.64153 48.353264 29.55491 49.794094 29.48151 51.23403 29.422285 52.672993 29.37881 54.1108 29.352652 55.547634 29.345558 56.983322 29.359749 57.605072 29.373585 57.61804 29.221487 57.836437 26.173342 58.010845 21.597244 58.017952 18.693539 57.946934 16.081406 57.844383 14.189138 57.696827 12.322918 57.54737 10.86875 57.35628 9.345355 57.17142 8.093174 56.95828 6.829593 56.937805 6.7161946 56.710182 5.5312023 56.41659 4.1687655 56.12184 2.942724 55.726597 1.4660592 55.310673 0.06907043 54.71953 -1.7121664 54.050846 -3.5155425 53.001633 -6.02846 51.629116 -8.914773 50.47874 -11.085491 50.47874 -11.085491" ;
            		:objectType = "gml:LinearRing" ;
            } // group gml\:exterior
          } // group gml\:surfaceMembers
        } // group eop\:multiExtentOf
      } // group om\:featureOfInterest

    group: eop\:metaDataProperty {

      // group attributes:
      		:objectType = "eop:EarthObservationMetaData" ;
      		:eop\:acquisitionType = "NOMINAL" ;
      		:eop\:identifier = "S5P_NRTI_L2__O3_____20240818T120300_20240818T120800_35484_03_020601_20240818T124850" ;
      		:eop\:doi = "N/A" ;
      		:eop\:parentIdentifier = "urn:ogc:def:EOP:ESA:SENTINEL.S5P_TROP_L2__O3____" ;
      		:eop\:productType = "S5P_NRTI_O3____" ;
      		:eop\:status = "ACQUIRED" ;
      		:eop\:productQualityStatus = "NOMINAL" ;
      		:eop\:productQualityDegradationTag = "NOT APPLICABLE" ;

      group: eop\:processing {

        // group attributes:
        		:objectType = "eop:ProcessingInformation" ;
        		:eop\:processingCenter = "PDGS-OP" ;
        		:eop\:processingDate = "2024-08-18" ;
        		:eop\:processingLevel = "L2" ;
        		:eop\:processorName = "upas-l2" ;
        		:eop\:processorVersion = "02.06.01" ;
        		:eop\:nativeProductFormat = "netCDF-4" ;
        		:eop\:processingMode = "NRTI" ;
        } // group eop\:processing
      } // group eop\:metaDataProperty
    } // group EOP_METADATA

  group: ISO_METADATA {

    // group attributes:
    		:gmd\:dateStamp = "2015-10-16" ;
    		:gmd\:fileIdentifier = "urn:ogc:def:EOP:ESA:SENTINEL.S5P_TROP_L2__O3____" ;
    		:gmd\:hierarchyLevelName = "EO Product Collection" ;
    		:gmd\:metadataStandardName = "ISO 19115-2 Geographic Information - Metadata Part 2 Extensions for imagery and gridded data" ;
    		:gmd\:metadataStandardVersion = "ISO 19115-2:2009(E), S5P profile" ;
    		:objectType = "gmi:MI_Metadata" ;

    group: gmd\:contact {

      // group attributes:
      		:gmd\:organisationName = "Copernicus Space Component Data Access System,  ESA, Services Coordinated Interface" ;
      		:objectType = "gmd:CI_ResponsibleParty" ;

      group: gmd\:role {

        // group attributes:
        		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_RoleCode" ;
        		:codeListValue = "pointOfContact" ;
        		:objectType = "gmd:CI_RoleCode" ;
        } // group gmd\:role

      group: gmd\:contactInfo {

        // group attributes:
        		:objectType = "gmd:CI_Contact" ;

        group: gmd\:address {

          // group attributes:
          		:gmd\:electronicMailAddress = "EOSupport@copernicus.esa.int" ;
          		:objectType = "gmd:CI_Address" ;
          } // group gmd\:address
        } // group gmd\:contactInfo
      } // group gmd\:contact

    group: gmd\:language {

      // group attributes:
      		:codeList = "http://www.loc.gov/standards/iso639-2/" ;
      		:codeListValue = "eng" ;
      		:objectType = "gmd:LanguageCode" ;
      } // group gmd\:language

    group: gmd\:characterSet {

      // group attributes:
      		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_CharacterSetCode" ;
      		:codeListValue = "utf8" ;
      		:objectType = "gmd:MD_CharacterSetCode" ;
      } // group gmd\:characterSet

    group: gmd\:hierarchyLevel {

      // group attributes:
      		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_ScopeCode" ;
      		:codeListValue = "series" ;
      		:objectType = "gmd:MD_ScopeCode" ;
      } // group gmd\:hierarchyLevel

    group: gmd\:dataQualityInfo {

      // group attributes:
      		:objectType = "gmd:DQ_DataQuality" ;

      group: gmd\:scope {

        // group attributes:
        		:objectType = "gmd:DQ_Scope" ;

        group: gmd\:level {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_ScopeCode" ;
          		:codeListValue = "dataset" ;
          		:objectType = "gmd:MD_ScopeCode" ;
          } // group gmd\:level
        } // group gmd\:scope

      group: gmd\:report {

        // group attributes:
        		:objectType = "gmd:DQ_DomainConsistency" ;

        group: gmd\:result {

          // group attributes:
          		:objectType = "gmd:DQ_ConformanceResult" ;
          		:gmd\:pass = "true" ;
          		:gmd\:explanation = "INSPIRE Data specification for orthoimagery is not yet officially published so conformity has not yet been evaluated" ;

          group: gmd\:specification {

            // group attributes:
            		:objectType = "gmd:CI_Citation" ;
            		:gmd\:title = "INSPIRE Data Specification on Orthoimagery - Guidelines, version 3.0rc3" ;

            group: gmd\:date {

              // group attributes:
              		:gmd\:date = "2013-02-04" ;
              		:objectType = "gmd:CI_Date" ;

              group: gmd\:dateType {

                // group attributes:
                		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                		:codeListValue = "publication" ;
                		:objectType = "gmd:CI_DateTypeCode" ;
                } // group gmd\:dateType
              } // group gmd\:date
            } // group gmd\:specification
          } // group gmd\:result
        } // group gmd\:report

      group: gmd\:lineage {

        // group attributes:
        		:objectType = "gmd:LI_Lineage" ;
        		:gmd\:statement = "L2 O3____ dataset produced by PDGS-OP from the S5P/TROPOMI L1B product" ;

        group: gmd\:processStep {

          // group attributes:
          		:objectType = "gmi:LE_ProcessStep" ;
          		:gmd\:description = "Processing of L1b to L2 O3____ data for orbit 35484 using the DLR-IMF processor version 02.06.01" ;

          group: gmi\:output {

            // group attributes:
            		:gmd\:description = "" ;
            		:objectType = "gmi:LE_Source" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L2" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:gmd\:title = "S5P_NRTI_L2__O3_____20240818T120300_20240818T120800_35484_03_020601_20240818T124850" ;
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "" ;
                		:objectType = "gmd:CI_DateTime" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:identifier {

                // group attributes:
                		:gmd\:code = "L2__O3____" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmd\:identifier
              } // group gmd\:sourceCitation
            } // group gmi\:output

          group: gmi\:report {

            // group attributes:
            		:gmi\:description = "Sentinel 5-precursor TROPOMI L1b processed to L2 data using the DLR-IMF L2 O3____ processor" ;
            		:gmi\:fileType = "netCDF-4" ;
            		:gmi\:name = "S5P_NRTI_L2__O3_____20240818T120300_20240818T120800_35484_03_020601_20240818T124850.nc" ;
            		:objectType = "gmi:LE_ProcessStepReport" ;
            } // group gmi\:report

          group: gmd\:source\#1 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_IR_UVN irradiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-08-18T12:49:05Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeList = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_IR_UVN irradiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_OFFL_L1B_IR_UVN_20240817T162923_20240817T181053_35473_03_020100_20240818T030032.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#1

          group: gmd\:source\#2 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_RA_BD1 radiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-08-18T12:49:05Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeList = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_RA_BD1 radiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD1_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#2

          group: gmd\:source\#3 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_RA_BD2 radiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-08-18T12:49:05Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeList = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_RA_BD2 radiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD2_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#3

          group: gmd\:source\#4 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_RA_BD3 radiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-08-18T12:49:05Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeList = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_RA_BD3 radiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD3_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#4

          group: gmd\:source\#5 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_RA_BD4 radiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-08-18T12:49:05Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeList = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_RA_BD4 radiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD4_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#5

          group: gmd\:source\#6 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_RA_BD5 radiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-08-18T12:49:05Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeList = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_RA_BD5 radiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD5_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#6

          group: gmd\:source\#7 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_RA_BD6 radiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-08-18T12:49:05Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeList = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_RA_BD6 radiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD6_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#7

          group: gmd\:source\#8 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_RA_BD7 radiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-08-18T12:49:05Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeList = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_RA_BD7 radiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD7_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#8

          group: gmd\:source\#9 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L1B L1B_RA_BD8 radiance product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L1B" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-08-18T12:49:05Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeList = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L1B L1B_RA_BD8 radiance product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD8_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#9

          group: gmd\:source\#10 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "TROPOMI L2 L2__CLOUD_ product" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "L2" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-08-18T12:49:05Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeList = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "TROPOMI L2 L2__CLOUD_ product" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_NRTI_L2__CLOUD__20240818T120300_20240818T120800_35484_03_020601_20240818T124206.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#10

          group: gmd\:source\#11 {

            // group attributes:
            		:objectType = "gmi:LE_Source" ;
            		:gmd\:description = "Auxiliary data" ;

            group: gmi\:processedLevel {

              // group attributes:
              		:gmd\:code = "N/A" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:processedLevel

            group: gmd\:sourceCitation {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2024-08-18T12:49:05Z" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeList = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date

              group: gmd\:title {

                // group attributes:
                		:gco\:characterString = "Auxiliary data" ;
                } // group gmd\:title

              group: gmd\:alternateTitle\#1 {

                // group attributes:
                		:gmx\:FileName = "S5P_NRTI_AUX_BGO3___20240815T205808_20240817T000320_20240818T000018.nc" ;
                } // group gmd\:alternateTitle\#1
              } // group gmd\:sourceCitation
            } // group gmd\:source\#11

          group: gmi\:processingInformation {

            // group attributes:
            		:objectType = "gmi:LE_Processing" ;

            group: gmi\:identifier {

              // group attributes:
              		:gmd\:code = "DLR-IMF L2 O3____ processor, version 02.06.01" ;
              		:objectType = "gmd:MD_Identifier" ;
              } // group gmi\:identifier

            group: gmi\:documentation\#1 {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;
              		:gmd\:title = "Sentinel-5 precursor/TROPOMI Ozone Total Column ATBD; S5P-L2-DLR-ATBD-400A; Release 1.0" ;
              		:doi = "N/A" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2016-02-01" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "publication" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date
              } // group gmi\:documentation\#1

            group: gmi\:documentation\#2 {

              // group attributes:
              		:objectType = "gmd:CI_Citation" ;
              		:gmd\:title = "Sentinel-5 precursor/TROPOMI Level 2 Product User Manual Ozone Total Column; S5P-L2-DLR-PUM-400A; Release 00.11.04" ;
              		:doi = "N/A" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2018-07-30" ;
                		:objectType = "gmd:CI_Date" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "publication" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date
              } // group gmi\:documentation\#2

            group: gmi\:softwareReference {

              // group attributes:
              		:gmd\:title = "UPAS L2 O3____ processor" ;
              		:objectType = "gmd:CI_Citation" ;

              group: gmd\:date {

                // group attributes:
                		:gmd\:date = "2023-11-10T14:17:48Z" ;
                		:objectType = "gmd:CI_DateTime" ;

                group: gmd\:dateType {

                  // group attributes:
                  		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                  		:codeListValue = "creation" ;
                  		:objectType = "gmd:CI_DateTypeCode" ;
                  } // group gmd\:dateType
                } // group gmd\:date
              } // group gmi\:softwareReference
            } // group gmi\:processingInformation
          } // group gmd\:processStep
        } // group gmd\:lineage
      } // group gmd\:dataQualityInfo

    group: gmd\:identificationInfo {

      // group attributes:
      		:gmd\:abstract = "" ;
      		:gmd\:credit = "The Sentinel 5 Precursor TROPOMI Level 2 products are developed with funding from the European Space Agency (ESA), the Netherlands Space Office (NSO), the Belgian Science Policy Office, the German Aerospace Center (DLR) and the Bayerisches Staatsministerium für Wirtschaft und Medien, Energie und Technologie (StMWi)." ;
      		:gmd\:language = "eng" ;
      		:gmd\:topicCategory = "climatologyMeteorologyAtmosphere" ;
      		:objectType = "gmd:MD_DataIdentification" ;

      group: gmd\:extent {

        // group attributes:
        		:objectType = "gmd:EX_Extent" ;

        group: gmd\:temporalElement {

          // group attributes:
          		:objectType = "gmd:EX_TemporalExtent" ;

          group: gmd\:extent {

            // group attributes:
            		:gml\:beginPosition = "2024-08-18T12:02:54Z" ;
            		:gml\:endPosition = "2024-08-18T12:08:07Z" ;
            		:objectType = "gml:TimePeriod" ;
            } // group gmd\:extent
          } // group gmd\:temporalElement

        group: gmd\:geographicElement {

          // group attributes:
          		:gmd\:eastBoundLongitude = 180.f ;
          		:gmd\:northBoundLatitude = 90.f ;
          		:gmd\:southBoundLatitude = -90.f ;
          		:gmd\:westBoundLongitude = -180.f ;
          		:gmd\:extentTypeCode = "true" ;
          		:objectType = "gmd:EX_GeographicBoundingBox" ;
          } // group gmd\:geographicElement
        } // group gmd\:extent

      group: gmd\:citation {

        // group attributes:
        		:gmd\:title = "" ;
        		:objectType = "gmd:CI_Citation" ;

        group: gmd\:date {

          // group attributes:
          		:gmd\:date = "2023-11-10T14:17:48Z" ;
          		:objectType = "gmd:CI_Date" ;

          group: gmd\:dateType {

            // group attributes:
            		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
            		:codeListValue = "creation" ;
            		:objectType = "gmd:CI_DateTypeCode" ;
            } // group gmd\:dateType
          } // group gmd\:date

        group: gmd\:identifier {

          // group attributes:
          		:gmd\:code = "urn:ogc:def:EOP:ESA:SENTINEL.S5P_TROP_L2__O3____" ;
          		:objectType = "gmd:MD_Identifier" ;
          } // group gmd\:identifier
        } // group gmd\:citation

      group: gmd\:characterSet {

        // group attributes:
        		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_CharacterSetCode" ;
        		:codeListValue = "utf8" ;
        		:objectType = "gmd:MD_CharacterSetCode" ;
        } // group gmd\:characterSet

      group: gmd\:pointOfContact {

        // group attributes:
        		:gmd\:organisationName = "Copernicus Space Component Data Access System,  ESA, Services Coordinated Interface" ;
        		:objectType = "gmd:CI_ResponsibleParty" ;

        group: gmd\:role {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_RoleCode" ;
          		:codeListValue = "distributor" ;
          		:objectType = "gmd:CI_RoleCode" ;
          } // group gmd\:role

        group: gmd\:contactInfo {

          // group attributes:
          		:objectType = "gmd:CI_Contact" ;

          group: gmd\:address {

            // group attributes:
            		:gmd\:electronicMailAddress = "EOSupport@copernicus.esa.int" ;
            		:objectType = "gmd:CI_Address" ;
            } // group gmd\:address
          } // group gmd\:contactInfo
        } // group gmd\:pointOfContact

      group: gmd\:spatialResolution {

        // group attributes:
        		:gmd\:distance = 7.f ;
        		:uom = "km" ;
        		:objectType = "gmd:MD_Resolution" ;
        } // group gmd\:spatialResolution

      group: gmd\:resourceConstraints {

        // group attributes:
        		:gmd\:useLimitation = "no conditions apply" ;
        		:objectType = "gmd:MD_LegalConstraints" ;

        group: gmd\:accessConstraints {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_RestrictionCode" ;
          		:codeListValue = "copyright" ;
          		:objectType = "gmd:MD_RestrictionCode" ;
          } // group gmd\:accessConstraints
        } // group gmd\:resourceConstraints

      group: gmd\:descriptiveKeywords\#2 {

        // group attributes:
        		:gmd\:keyword\#1 = "" ;
        		:objectType = "gmd:MD_Keywords" ;

        group: gmd\:thesaurusName {

          // group attributes:
          		:gmd\:title = "CF Standard Name Table v29" ;
          		:xlink\:href = "http://cfconventions.org/standard-names.html" ;
          		:objectType = "gmd:CI_Citation" ;

          group: gmd\:date {

            // group attributes:
            		:gmd\:date = "2015-07-08" ;
            		:objectType = "gmd:CI_Date" ;

            group: gmd\:dateType {

              // group attributes:
              		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
              		:codeListValue = "publication" ;
              		:objectType = "gmd:CI_DateTypeCode" ;
              } // group gmd\:dateType
            } // group gmd\:date
          } // group gmd\:thesaurusName
        } // group gmd\:descriptiveKeywords\#2

      group: gmd\:descriptiveKeywords\#1 {

        // group attributes:
        		:gmd\:keyword\#1 = "Atmospheric conditions" ;
        		:objectType = "gmd:MD_Keywords" ;

        group: gmd\:type {

          // group attributes:
          		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_KeywordTypeCode" ;
          		:codeListValue = "theme" ;
          		:objectType = "gmd:MD_KeywordTypeCode" ;
          } // group gmd\:type

        group: gmd\:thesaurusName {

          // group attributes:
          		:gmd\:title = "GEMET - INSPIRE themes, version 1.0" ;
          		:objectType = "gmd:CI_Citation" ;

          group: gmd\:date {

            // group attributes:
            		:gmd\:date = "2008-06-01" ;
            		:objectType = "gmd:CI_Date" ;

            group: gmd\:dateType {

              // group attributes:
              		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
              		:codeListValue = "publication" ;
              		:objectType = "gmd:CI_DateTypeCode" ;
              } // group gmd\:dateType
            } // group gmd\:date
          } // group gmd\:thesaurusName
        } // group gmd\:descriptiveKeywords\#1

      group: gmd\:spatialRepresentationType {

        // group attributes:
        		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#MD_SpatialRepresentationTypeCode" ;
        		:codeListValue = "grid" ;
        		:objectType = "gmd:MD_SpatialRepresentationTypeCode" ;
        } // group gmd\:spatialRepresentationType
      } // group gmd\:identificationInfo

    group: gmi\:acquisitionInformation {

      // group attributes:
      		:objectType = "gmi:MI_AcquisitionInformation" ;

      group: gmi\:platform {

        // group attributes:
        		:gmi\:description = "Sentinel 5 Precursor" ;
        		:objectType = "gmi:MI_Platform" ;

        group: gmi\:instrument {

          // group attributes:
          		:objectType = "gmi:MI_Instrument" ;
          		:gmi\:type = "UV-VIS-NIR-SWIR imaging spectrometer" ;

          group: gmi\:identifier {

            // group attributes:
            		:gmd\:code = "TROPOMI" ;
            		:gmd\:codeSpace = "http://www.esa.int/" ;
            		:objectType = "gmd:RS_Identifier" ;
            } // group gmi\:identifier
          } // group gmi\:instrument

        group: gmi\:identifier {

          // group attributes:
          		:gmd\:code = "S5P" ;
          		:gmd\:codeSpace = "http://www.esa.int/" ;
          		:objectType = "gmd:RS_Identifier" ;
          } // group gmi\:identifier
        } // group gmi\:platform
      } // group gmi\:acquisitionInformation
    } // group ISO_METADATA

  group: QA_STATISTICS {
    dimensions:
    	vertices = 2 ;
    	histogram_axis = 100 ;
    	pdf_axis = 400 ;
    variables:
    	float histogram_axis(histogram_axis) ;
    		histogram_axis:_FillValue = 9.96921e+36f ;
    		histogram_axis:units = "1" ;
    		histogram_axis:bounds = "histogram_bounds" ;
    	float pdf_axis(pdf_axis) ;
    		pdf_axis:_FillValue = 9.96921e+36f ;
    		pdf_axis:units = "1" ;
    		pdf_axis:bounds = "pdf_bounds" ;
    	int ozone_total_column_histogram(histogram_axis) ;
    		ozone_total_column_histogram:_FillValue = -2147483647 ;
    		ozone_total_column_histogram:comment = "Histogram of the total column O3 in the current granule" ;
    	float ozone_total_column_pdf(pdf_axis) ;
    		ozone_total_column_pdf:_FillValue = 9.96921e+36f ;
    		ozone_total_column_pdf:comment = "Probability density function of the total column O3 in the current granule" ;
    	int vertices(vertices) ;
    		vertices:units = "1" ;
    		vertices:long_name = "vertices dimension index" ;

    // group attributes:
    		:number_of_groundpixels = 160650 ;
    		:number_of_processed_pixels = 160650 ;
    		:number_of_successfully_processed_pixels = 160293 ;
    		:number_of_rejected_pixels_not_enough_spectrum = 0 ;
    		:number_of_failed_retrievals = 0 ;
    		:number_of_ground_pixels_with_warnings = 0 ;
    		:number_of_radiance_missing_occurrences = 0 ;
    		:number_of_irradiance_missing_occurrences = 0 ;
    		:number_of_input_spectrum_missing_occurrences = 0 ;
    		:number_of_reflectance_range_error_occurrences = 0 ;
    		:number_of_ler_range_error_occurrences = 0 ;
    		:number_of_snr_range_error_occurrences = 0 ;
    		:number_of_sza_range_error_occurrences = 0 ;
    		:number_of_vza_range_error_occurrences = 0 ;
    		:number_of_lut_range_error_occurrences = 0 ;
    		:number_of_ozone_range_error_occurrences = 0 ;
    		:number_of_wavelength_offset_error_occurrences = 0 ;
    		:number_of_initialization_error_occurrences = 0 ;
    		:number_of_memory_error_occurrences = 0 ;
    		:number_of_assertion_error_occurrences = 0 ;
    		:number_of_io_error_occurrences = 0 ;
    		:number_of_numerical_error_occurrences = 0 ;
    		:number_of_lut_error_occurrences = 0 ;
    		:number_of_ISRF_error_occurrences = 0 ;
    		:number_of_convergence_error_occurrences = 0 ;
    		:number_of_cloud_filter_convergence_error_occurrences = 0 ;
    		:number_of_max_iteration_convergence_error_occurrences = 0 ;
    		:number_of_aot_lower_boundary_convergence_error_occurrences = 0 ;
    		:number_of_other_boundary_convergence_error_occurrences = 0 ;
    		:number_of_geolocation_error_occurrences = 0 ;
    		:number_of_ch4_noscat_zero_error_occurrences = 0 ;
    		:number_of_h2o_noscat_zero_error_occurrences = 0 ;
    		:number_of_max_optical_thickness_error_occurrences = 0 ;
    		:number_of_aerosol_boundary_error_occurrences = 0 ;
    		:number_of_boundary_hit_error_occurrences = 0 ;
    		:number_of_chi2_error_occurrences = 0 ;
    		:number_of_svd_error_occurrences = 0 ;
    		:number_of_dfs_error_occurrences = 0 ;
    		:number_of_radiative_transfer_error_occurrences = 0 ;
    		:number_of_optimal_estimation_error_occurrences = 0 ;
    		:number_of_profile_error_occurrences = 0 ;
    		:number_of_cloud_error_occurrences = 0 ;
    		:number_of_model_error_occurrences = 0 ;
    		:number_of_number_of_input_data_points_too_low_error_occurrences = 0 ;
    		:number_of_cloud_pressure_spread_too_low_error_occurrences = 0 ;
    		:number_of_cloud_too_low_level_error_occurrences = 0 ;
    		:number_of_generic_range_error_occurrences = 0 ;
    		:number_of_generic_exception_occurrences = 357 ;
    		:number_of_input_spectrum_alignment_error_occurrences = 0 ;
    		:number_of_abort_error_occurrences = 0 ;
    		:number_of_wrong_input_type_error_occurrences = 0 ;
    		:number_of_wavelength_calibration_error_occurrences = 0 ;
    		:number_of_coregistration_error_occurrences = 0 ;
    		:number_of_slant_column_density_error_occurrences = 0 ;
    		:number_of_airmass_factor_error_occurrences = 0 ;
    		:number_of_vertical_column_density_error_occurrences = 0 ;
    		:number_of_signal_to_noise_ratio_error_occurrences = 0 ;
    		:number_of_configuration_error_occurrences = 0 ;
    		:number_of_key_error_occurrences = 0 ;
    		:number_of_saturation_error_occurrences = 0 ;
    		:number_of_solar_eclipse_filter_occurrences = 0 ;
    		:number_of_cloud_filter_occurrences = 0 ;
    		:number_of_altitude_consistency_filter_occurrences = 0 ;
    		:number_of_altitude_roughness_filter_occurrences = 0 ;
    		:number_of_sun_glint_filter_occurrences = 0 ;
    		:number_of_mixed_surface_type_filter_occurrences = 0 ;
    		:number_of_snow_ice_filter_occurrences = 0 ;
    		:number_of_aai_filter_occurrences = 0 ;
    		:number_of_cloud_fraction_fresco_filter_occurrences = 0 ;
    		:number_of_aai_scene_albedo_filter_occurrences = 0 ;
    		:number_of_small_pixel_radiance_std_filter_occurrences = 0 ;
    		:number_of_cloud_fraction_viirs_filter_occurrences = 0 ;
    		:number_of_cirrus_reflectance_viirs_filter_occurrences = 0 ;
    		:number_of_cf_viirs_swir_ifov_filter_occurrences = 0 ;
    		:number_of_cf_viirs_swir_ofova_filter_occurrences = 0 ;
    		:number_of_cf_viirs_swir_ofovb_filter_occurrences = 0 ;
    		:number_of_cf_viirs_swir_ofovc_filter_occurrences = 0 ;
    		:number_of_cf_viirs_nir_ifov_filter_occurrences = 0 ;
    		:number_of_cf_viirs_nir_ofova_filter_occurrences = 0 ;
    		:number_of_cf_viirs_nir_ofovb_filter_occurrences = 0 ;
    		:number_of_cf_viirs_nir_ofovc_filter_occurrences = 0 ;
    		:number_of_refl_cirrus_viirs_swir_filter_occurrences = 0 ;
    		:number_of_refl_cirrus_viirs_nir_filter_occurrences = 0 ;
    		:number_of_diff_refl_cirrus_viirs_filter_occurrences = 0 ;
    		:number_of_ch4_noscat_ratio_filter_occurrences = 0 ;
    		:number_of_ch4_noscat_ratio_std_filter_occurrences = 0 ;
    		:number_of_h2o_noscat_ratio_filter_occurrences = 0 ;
    		:number_of_h2o_noscat_ratio_std_filter_occurrences = 0 ;
    		:number_of_diff_psurf_fresco_ecmwf_filter_occurrences = 0 ;
    		:number_of_psurf_fresco_stdv_filter_occurrences = 0 ;
    		:number_of_ocean_filter_occurrences = 0 ;
    		:number_of_time_range_filter_occurrences = 0 ;
    		:number_of_pixel_or_scanline_index_filter_occurrences = 0 ;
    		:number_of_geographic_region_filter_occurrences = 0 ;
    		:number_of_input_spectrum_warning_occurrences = 0 ;
    		:number_of_wavelength_calibration_warning_occurrences = 0 ;
    		:number_of_extrapolation_warning_occurrences = 0 ;
    		:number_of_sun_glint_warning_occurrences = 0 ;
    		:number_of_south_atlantic_anomaly_warning_occurrences = 0 ;
    		:number_of_sun_glint_correction_occurrences = 0 ;
    		:number_of_snow_ice_warning_occurrences = 0 ;
    		:number_of_cloud_warning_occurrences = 53699 ;
    		:number_of_AAI_warning_occurrences = 0 ;
    		:number_of_pixel_level_input_data_missing_occurrences = 0 ;
    		:number_of_data_range_warning_occurrences = 0 ;
    		:number_of_low_cloud_fraction_warning_occurrences = 0 ;
    		:number_of_altitude_consistency_warning_occurrences = 0 ;
    		:number_of_signal_to_noise_ratio_warning_occurrences = 0 ;
    		:number_of_deconvolution_warning_occurrences = 0 ;
    		:number_of_so2_volcanic_origin_likely_warning_occurrences = 0 ;
    		:number_of_so2_volcanic_origin_certain_warning_occurrences = 0 ;
    		:number_of_interpolation_warning_occurrences = 0 ;
    		:number_of_saturation_warning_occurrences = 0 ;
    		:number_of_high_sza_warning_occurrences = 0 ;
    		:number_of_cloud_retrieval_warning_occurrences = 1430 ;
    		:number_of_cloud_inhomogeneity_warning_occurrences = 33525 ;
    		:global_processing_warnings = "None" ;
    		:time_for_algorithm_initialization = 2.38 ;
    		:time_for_processing = 33.04 ;
    		:time_per_pixel = 0.000206 ;
    		:time_standard_deviation_per_pixel = 0.000206 ;
    } // group QA_STATISTICS

  group: GRANULE_DESCRIPTION {

    // group attributes:
    		:GranuleStart = "2024-08-18T12:02:54Z" ;
    		:GranuleEnd = "2024-08-18T12:08:07Z" ;
    		:InstrumentName = "TROPOMI" ;
    		:MissionName = "Sentinel-5 precursor" ;
    		:MissionShortName = "S5P" ;
    		:ProcessLevel = "2" ;
    		:ProcessingCenter = "PDGS-OP" ;
    		:ProcessingNode = "s5p-ops2-nrt-pn05" ;
    		:ProcessorVersion = "02.06.01" ;
    		:ProductFormatVersion = 1 ;
    		:ProcessingMode = "Near-realtime" ;
    		:CollectionIdentifier = "" ;
    		:ProductShortName = "L2__O3____" ;
    } // group GRANULE_DESCRIPTION

  group: ESA_METADATA {

    group: earth_explorer_header {

      // group attributes:
      		:objectType = "Earth_Explorer_Header" ;

      group: fixed_header {

        // group attributes:
        		:objectType = "Fixed_Header" ;
        		:File_Name = "S5P_NRTI_L2__O3_____20240818T120300_20240818T120800_35484_03_020601_20240818T124850" ;
        		:File_Description = "" ;
        		:Notes = "" ;
        		:Mission = "S5P" ;
        		:File_Class = "NRTI" ;
        		:File_Type = "L2__O3____" ;
        		:File_Version = 0 ;

        group: source {

          // group attributes:
          		:objectType = "Source" ;
          		:System = "PDGS-OP" ;
          		:Creator = "upas-l2" ;
          		:Creator_Version = "02.06.01" ;
          		:Creation_Date = "UTC=2024-08-18T12:49:05" ;
          } // group source

        group: validity_period {

          // group attributes:
          		:objectType = "Validity_Period" ;
          		:Validity_Start = "UTC=2024-08-18T12:02:54" ;
          		:Validity_Stop = "UTC=2024-08-18T12:08:07" ;
          } // group validity_period
        } // group fixed_header

      group: variable_header {

        // group attributes:
        		:objectType = "Variable_Header" ;

        group: gmd\:lineage {

          // group attributes:
          		:objectType = "gmd:LI_Lineage" ;
          		:gmd\:statement = "L2 O3____ dataset produced by PDGS-OP from the S5P/TROPOMI L1B product" ;

          group: gmd\:processStep {

            // group attributes:
            		:objectType = "gmi:LE_ProcessStep" ;
            		:gmd\:description = "Processing of L1b to L2 O3____ data for orbit 35484 using the DLR-IMF processor version 02.06.01" ;

            group: gmi\:output {

              // group attributes:
              		:gmd\:description = "" ;
              		:objectType = "gmi:LE_Source" ;

              group: gmd\:sourceCitation {

                // group attributes:
                		:gmd\:title = "S5P_NRTI_L2__O3_____20240818T120300_20240818T120800_35484_03_020601_20240818T124850" ;
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "" ;
                  		:objectType = "gmd:CI_DateTime" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:identifier {

                  // group attributes:
                  		:gmd\:code = "L2__O3____" ;
                  		:objectType = "gmd:MD_Identifier" ;
                  } // group gmd\:identifier
                } // group gmd\:sourceCitation

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L2" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel
              } // group gmi\:output

            group: gmi\:report {

              // group attributes:
              		:gmi\:description = "Sentinel 5-precursor TROPOMI L1b processed to L2 data using the DLR-IMF L2 O3____ processor" ;
              		:gmi\:fileType = "netCDF-4" ;
              		:gmi\:name = "S5P_NRTI_L2__O3_____20240818T120300_20240818T120800_35484_03_020601_20240818T124850.nc" ;
              		:objectType = "gmi:LE_ProcessStepReport" ;
              } // group gmi\:report

            group: gmd\:source\#1 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_IR_UVN irradiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-08-18T12:49:05Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeList = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_IR_UVN irradiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_OFFL_L1B_IR_UVN_20240817T162923_20240817T181053_35473_03_020100_20240818T030032.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#1

            group: gmd\:source\#2 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_RA_BD1 radiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-08-18T12:49:05Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeList = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_RA_BD1 radiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD1_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#2

            group: gmd\:source\#3 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_RA_BD2 radiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-08-18T12:49:05Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeList = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_RA_BD2 radiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD2_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#3

            group: gmd\:source\#4 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_RA_BD3 radiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-08-18T12:49:05Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeList = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_RA_BD3 radiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD3_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#4

            group: gmd\:source\#5 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_RA_BD4 radiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-08-18T12:49:05Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeList = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_RA_BD4 radiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD4_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#5

            group: gmd\:source\#6 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_RA_BD5 radiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-08-18T12:49:05Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeList = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_RA_BD5 radiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD5_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#6

            group: gmd\:source\#7 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_RA_BD6 radiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-08-18T12:49:05Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeList = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_RA_BD6 radiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD6_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#7

            group: gmd\:source\#8 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_RA_BD7 radiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-08-18T12:49:05Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeList = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_RA_BD7 radiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD7_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#8

            group: gmd\:source\#9 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L1B L1B_RA_BD8 radiance product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L1B" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-08-18T12:49:05Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeList = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L1B L1B_RA_BD8 radiance product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_NRTI_L1B_RA_BD8_20240818T120254_20240818T120806_35484_03_020100_20240818T122756.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#9

            group: gmd\:source\#10 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "TROPOMI L2 L2__CLOUD_ product" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "L2" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-08-18T12:49:05Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeList = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "TROPOMI L2 L2__CLOUD_ product" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_NRTI_L2__CLOUD__20240818T120300_20240818T120800_35484_03_020601_20240818T124206.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#10

            group: gmd\:source\#11 {

              // group attributes:
              		:objectType = "gmi:LE_Source" ;
              		:gmd\:description = "Auxiliary data" ;

              group: gmi\:processedLevel {

                // group attributes:
                		:gmd\:code = "N/A" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:processedLevel

              group: gmd\:sourceCitation {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2024-08-18T12:49:05Z" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeListValue = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeList = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date

                group: gmd\:title {

                  // group attributes:
                  		:gco\:characterString = "Auxiliary data" ;
                  } // group gmd\:title

                group: gmd\:alternateTitle\#1 {

                  // group attributes:
                  		:gmx\:FileName = "S5P_NRTI_AUX_BGO3___20240815T205808_20240817T000320_20240818T000018.nc" ;
                  } // group gmd\:alternateTitle\#1
                } // group gmd\:sourceCitation
              } // group gmd\:source\#11

            group: gmi\:processingInformation {

              // group attributes:
              		:objectType = "gmi:LE_Processing" ;

              group: gmi\:identifier {

                // group attributes:
                		:gmd\:code = "DLR-IMF L2 O3____ processor, version 02.06.01" ;
                		:objectType = "gmd:MD_Identifier" ;
                } // group gmi\:identifier

              group: gmi\:documentation\#2 {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;
                		:gmd\:title = "Sentinel-5 precursor/TROPOMI Level 2 Product User Manual Ozone Total Column; S5P-L2-DLR-PUM-400A; Release 00.11.04" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2018-07-30" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "publication" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:documentation\#2

              group: gmi\:documentation\#1 {

                // group attributes:
                		:objectType = "gmd:CI_Citation" ;
                		:gmd\:title = "Sentinel-5 precursor/TROPOMI Ozone Total Column ATBD; S5P-L2-DLR-ATBD-400A; Release 1.0" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2016-02-01" ;
                  		:objectType = "gmd:CI_Date" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "publication" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:documentation\#1

              group: gmi\:softwareReference {

                // group attributes:
                		:gmd\:title = "UPAS L2 O3____ processor" ;
                		:objectType = "gmd:CI_Citation" ;

                group: gmd\:date {

                  // group attributes:
                  		:gmd\:date = "2023-11-10T14:17:48Z" ;
                  		:objectType = "gmd:CI_DateTime" ;

                  group: gmd\:dateType {

                    // group attributes:
                    		:codeList = "http://www.isotc211.org/2005/resources/Codelist/gmxCodelists.xml#CI_DateTypeCode" ;
                    		:codeListValue = "creation" ;
                    		:objectType = "gmd:CI_DateTypeCode" ;
                    } // group gmd\:dateType
                  } // group gmd\:date
                } // group gmi\:softwareReference
              } // group gmi\:processingInformation
            } // group gmd\:processStep
          } // group gmd\:lineage
        } // group variable_header
      } // group earth_explorer_header
    } // group ESA_METADATA
  } // group METADATA
}
